module RGB_led (
    input sys_clk,
    input sys_rst_n,
    input [7:0] in_R,
    input [7:0] in_G, 
    input [7:0] in_B,
    output R, G, B
);

PWM pwmR (
    .clk(sys_clk),
    .sys_rst_n(sys_rst_n),
    .duty_cycle(in_R),
    .out(R)
);
PWM pwmG (
    .clk(sys_clk),
    .sys_rst_n(sys_rst_n),
    .duty_cycle(in_G),
    .out(G)
);
PWM pwmB (
    .clk(sys_clk),
    .sys_rst_n(sys_rst_n),
    .duty_cycle(in_B),
    .out(B)
);

endmodule

module PWM (
    input clk,
    input sys_rst_n,
    input [7:0] duty_cycle, // 1 ~ 100
    output reg out
);

wire [6:0] cnt; // 1~100

always @(*) begin
    if (!sys_rst_n) begin
        out = 0;
    end else begin
        out = (cnt <= duty_cycle);
    end
end

PWM_counter #(
    .Max(100),
    .Min(1)
) PWM_cnt (
    .clk(clk),
    .enable(1'b1),
    .sys_rst_n(sys_rst_n),
    .U_D(1'b0), // 1: down, 0: up
    .cnt(cnt)
);

endmodule

module PWM_counter #(
    parameter Max = 15,
    parameter Min = 0
)(
    input clk,
    input enable,
    input sys_rst_n,
    input U_D, // 1: down, 0: up
    output reg [$clog2(Max + 1) - 1:0] cnt
);

    reg dir;

    always @(posedge clk or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            cnt <= Min;
        end else if (!enable) begin
            cnt <= cnt;
        end else if (cnt == Max && dir == 0) begin
            cnt <= Min;
        end else if (cnt == Min && dir == 1) begin
            cnt <= Max;
        end else begin
            cnt <= (dir) ? cnt - 1 : cnt + 1;
        end
    end

    always @(negedge clk or negedge sys_rst_n) begin
        if (!sys_rst_n) begin
            dir <= 1'b0;
        end else begin
            dir <= U_D;
        end
    end

endmodule
